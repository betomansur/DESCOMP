library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 4;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
		  
		  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant AND1 : std_logic_vector(3 downto 0) := "1011";

		  
		  
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:tmp(0) := x"5" & '1' & x"FF";   -- STA @511
tmp(0) := x"0" & '0' & x"00";   -- NOP
tmp(1) := x"4" & '0' & x"00";   -- LDI $0       # Carrega o valor 0 no acumulador
tmp(2) := x"5" & '1' & x"FE";   -- STA @510     # Limpa a leitura de KEY0 escrevendo no endereÃ§o de memÃ³ria 510
tmp(3) := x"5" & '1' & x"FF";   -- STA @511     # Limpa a leitura de KEY1 escrevendo no endereÃ§o de memÃ³ria 511
tmp(4) := x"5" & '1' & x"FD";   -- STA @509     # Limpa a leitura de FPGA_RESET escrevendo no endereÃ§o de memÃ³ria 509
tmp(5) := x"5" & '0' & x"00";   -- STA @0       # Define o valor no endereÃ§o de memÃ³ria 0 como 0
tmp(6) := x"5" & '1' & x"20";   -- STA @288     # Limpa o display HEX0
tmp(7) := x"5" & '1' & x"21";   -- STA @289     # Limpa o display HEX1
tmp(8) := x"5" & '1' & x"22";   -- STA @290     # Limpa o display HEX2
tmp(9) := x"5" & '1' & x"23";   -- STA @291     # Limpa o display HEX3
tmp(10) := x"5" & '1' & x"24";  -- STA @292     # Limpa o display HEX4
tmp(11) := x"5" & '1' & x"25";  -- STA @293     # Limpa o display HEX5
tmp(12) := x"5" & '1' & x"00";  -- STA @256     # Limpa todos os LEDs de LEDR0 a LEDR7
tmp(13) := x"5" & '1' & x"01";  -- STA @257     # Limpa LEDR8
tmp(14) := x"5" & '1' & x"02";  -- STA @258     # Limpa LEDR9
tmp(15) := x"5" & '1' & x"40";  -- STA @320     # Limpa o valor lido dos switches SW0 a SW7
tmp(16) := x"5" & '1' & x"41";  -- STA @321     # Limpa o valor lido do switch SW8
tmp(17) := x"5" & '1' & x"42";  -- STA @322     # Limpa o valor lido do switch SW9
tmp(18) := x"5" & '0' & x"10";  -- STA @16      # Reseta o contador no endereÃ§o de memÃ³ria para Unidade
tmp(19) := x"5" & '0' & x"11";  -- STA @17      # Reseta o contador no endereÃ§o de memÃ³ria para Dezenas
tmp(20) := x"5" & '0' & x"12";  -- STA @18      # Reseta o contador no endereÃ§o de memÃ³ria para Centenas
tmp(21) := x"5" & '0' & x"13";  -- STA @19      # Reseta o contador no endereÃ§o de memÃ³ria para Milhares
tmp(22) := x"5" & '0' & x"14";  -- STA @20      # Reseta o contador no endereÃ§o de memÃ³ria para Centenas de Milhar
tmp(23) := x"5" & '0' & x"15";  -- STA @21      # Reseta o contador no endereÃ§o de memÃ³ria para Dezenas de Milhar
tmp(24) := x"5" & '0' & x"20";  -- STA @32      # Reseta os limites de contagem para Unidade
tmp(25) := x"5" & '0' & x"21";  -- STA @33      # Reseta os limites de contagem para Dezenas
tmp(26) := x"5" & '0' & x"22";  -- STA @34      # Reseta os limites de contagem para Centenas
tmp(27) := x"5" & '0' & x"23";  -- STA @35      # Reseta os limites de contagem para Unidade de Milhar
tmp(28) := x"5" & '0' & x"24";  -- STA @36      # Reseta os limites de contagem para Dezenas de Milhar
tmp(29) := x"5" & '0' & x"25";  -- STA @37      # Reseta os limites de contagem para Centenas de Milhar
tmp(30) := x"5" & '0' & x"1B";  -- STA @27      # Limpa a flag de limite
tmp(31) := x"4" & '0' & x"01";  -- LDI $1       # Carrega o valor 1 no acumulador
tmp(32) := x"5" & '0' & x"01";  -- STA @1       # Define o valor no endereÃ§o de memÃ³ria 1 como 1
tmp(33) := x"4" & '0' & x"0A";  -- LDI $10      # Carrega o valor 10 no acumulador
tmp(34) := x"5" & '0' & x"0A";  -- STA @10      # Define o valor no endereÃ§o de memÃ³ria 10 como 10
tmp(35) := x"4" & '0' & x"0F";  -- LDI $15      # Carrega o valor 15 no acumulador
tmp(36) := x"5" & '0' & x"0F";  -- STA @15      # Define o valor no endereÃ§o de memÃ³ria 15 como 15
tmp(37) := x"0" & '0' & x"00"; -- NOP #LOOP:pra pular na linha 37
tmp(38) := x"1" & '1' & x"60";  -- LDA @352     # LÃª o estado da chave KEY0
tmp(39) := x"B" & '0' & x"01";  -- AND @1       # Aplica mÃ¡scara para isolar o bit 0
tmp(40) := x"8" & '0' & x"00";  -- CEQ @0       # Compara com 0, continua se KEY0 nÃ£o estiver pressionado
tmp(41) := x"7" & '0' & x"2C";  -- JEQ @PASSAKEY0       # Salta se igual, ou seja, KEY0 nÃ£o pressionado
tmp(42) := x"9" & '0' & x"3B";  -- JSR @INCREMENTA      # Chama sub-rotina para incrementar contadores
tmp(43) := x"9" & '1' & x"03";  -- JSR @VERIFICARLIMITE         # Chama sub-rotina para verificar se os contadores atingiram limites
tmp(44) := x"0" & '0' & x"00"; -- NOP #PASSAKEY0:pra pular na linha 44
tmp(45) := x"1" & '1' & x"61";  -- LDA @353     # LÃª o estado da chave KEY1
tmp(46) := x"B" & '0' & x"01";  -- AND @1       # Aplica mÃ¡scara para isolar o bit 0
tmp(47) := x"8" & '0' & x"00";  -- CEQ @0       # Compara com 0, continua se KEY1 nÃ£o estiver pressionado
tmp(48) := x"7" & '0' & x"32";  -- JEQ @PASSAKEY1       # Salta se igual, ou seja, KEY1 nÃ£o pressionado
tmp(49) := x"9" & '0' & x"91";  -- JSR @CONFIGURACAO    # Chama sub-rotina de configuraÃ§Ã£o se KEY1 estiver pressionado
tmp(50) := x"0" & '0' & x"00"; -- NOP #PASSAKEY1:pra pular na linha 50
tmp(51) := x"1" & '1' & x"64";  -- LDA @356     # LÃª o estado do botÃ£o FPGA_RESET
tmp(52) := x"B" & '0' & x"01";  -- AND @1       # Aplica mÃ¡scara para isolar o bit 0
tmp(53) := x"8" & '0' & x"00";  -- CEQ @0       # Compara com 0, continua se FPGA_RESET nÃ£o estiver pressionado
tmp(54) := x"7" & '0' & x"38";  -- JEQ @PASSAFPGARESET  # Salta se igual, ou seja, FPGA_RESET nÃ£o pressionado
tmp(55) := x"9" & '0' & x"F0";  -- JSR @REINICIACONTAGEM        # Chama sub-rotina para reiniciar a contagem
tmp(56) := x"0" & '0' & x"00"; -- NOP #PASSAFPGARESET:pra pular na linha 56
tmp(57) := x"6" & '0' & x"25";  -- JMP @LOOP    # Volta ao inÃ­cio do loop principal
tmp(58) := x"0" & '0' & x"00";  -- NOP
tmp(59) := x"0" & '0' & x"00"; -- NOP #INCREMENTA:pra pular na linha 59
tmp(60) := x"5" & '1' & x"FF";  -- STA @511     # Limpa a leitura de KEY0
tmp(61) := x"1" & '0' & x"1B";  -- LDA @27      # Carrega a flag de limite
tmp(62) := x"8" & '0' & x"01";  -- CEQ @1       # Compara com 1
tmp(63) := x"7" & '0' & x"8F";  -- JEQ @RETORNOINCREMENTA       # Salta se igual, ou seja, hÃ¡ limite alcanÃ§ado
tmp(64) := x"0" & '0' & x"00";  -- NOP
tmp(65) := x"1" & '0' & x"10";  -- LDA @16      # Carrega valor da Unidade
tmp(66) := x"2" & '0' & x"01";  -- SOMA @1      # Soma 1
tmp(67) := x"5" & '0' & x"10";  -- STA @16      # Armazena o novo valor da Unidade
tmp(68) := x"1" & '0' & x"10";  -- LDA @16
tmp(69) := x"8" & '0' & x"0A";  -- CEQ @10      # Compara se a Unidade Ã© igual a 10
tmp(70) := x"7" & '0' & x"4A";  -- JEQ @INCREMENTADEZENA        # Salta se igual para incrementar a Dezena
tmp(71) := x"1" & '0' & x"10";  -- LDA @16
tmp(72) := x"5" & '1' & x"20";  -- STA @288     # Atualiza display HEX0
tmp(73) := x"6" & '0' & x"8F";  -- JMP @RETORNOINCREMENTA
tmp(74) := x"0" & '0' & x"00"; -- NOP #INCREMENTADEZENA:pra pular na linha 74
tmp(75) := x"1" & '0' & x"00";  -- LDA @0
tmp(76) := x"5" & '0' & x"10";  -- STA @16      # Reseta a Unidade
tmp(77) := x"5" & '1' & x"20";  -- STA @288     # Atualiza display HEX0
tmp(78) := x"1" & '0' & x"11";  -- LDA @17
tmp(79) := x"2" & '0' & x"01";  -- SOMA @1      # Soma 1 na Dezena
tmp(80) := x"5" & '0' & x"11";  -- STA @17      # Armazena o novo valor da Dezena
tmp(81) := x"1" & '0' & x"11";  -- LDA @17
tmp(82) := x"8" & '0' & x"0A";  -- CEQ @10      # Compara se a Dezena Ã© igual a 10
tmp(83) := x"7" & '0' & x"57";  -- JEQ @INCREMENTACENTENA       # Salta se igual para incrementar a Centena
tmp(84) := x"1" & '0' & x"11";  -- LDA @17
tmp(85) := x"5" & '1' & x"21";  -- STA @289     # Atualiza display HEX1
tmp(86) := x"6" & '0' & x"8F";  -- JMP @RETORNOINCREMENTA
tmp(87) := x"0" & '0' & x"00"; -- NOP #INCREMENTACENTENA:pra pular na linha 87
tmp(88) := x"1" & '0' & x"00";  -- LDA @0
tmp(89) := x"5" & '0' & x"11";  -- STA @17      # Reseta a Dezena
tmp(90) := x"5" & '1' & x"21";  -- STA @289     # Atualiza display HEX1
tmp(91) := x"1" & '0' & x"12";  -- LDA @18
tmp(92) := x"2" & '0' & x"01";  -- SOMA @1      # Soma 1 na Centena
tmp(93) := x"5" & '0' & x"12";  -- STA @18      # Armazena o novo valor da Centena
tmp(94) := x"1" & '0' & x"12";  -- LDA @18
tmp(95) := x"8" & '0' & x"0A";  -- CEQ @10      # Compara se a Centena Ã© igual a 10
tmp(96) := x"7" & '0' & x"64";  -- JEQ @INCREMENTAMILHAR        # Salta se igual para incrementar o Milhar
tmp(97) := x"1" & '0' & x"12";  -- LDA @18
tmp(98) := x"5" & '1' & x"22";  -- STA @290     # Atualiza display HEX2
tmp(99) := x"6" & '0' & x"8F";  -- JMP @RETORNOINCREMENTA
tmp(100) := x"0" & '0' & x"00"; -- NOP #INCREMENTAMILHAR:pra pular na linha 100
tmp(101) := x"1" & '0' & x"00"; -- LDA @0
tmp(102) := x"5" & '0' & x"12"; -- STA @18      # Reseta a Centena
tmp(103) := x"5" & '1' & x"22"; -- STA @290     # Atualiza display HEX2
tmp(104) := x"1" & '0' & x"13"; -- LDA @19
tmp(105) := x"2" & '0' & x"01"; -- SOMA @1      # Soma 1 no Milhar
tmp(106) := x"5" & '0' & x"13"; -- STA @19      # Armazena o novo valor do Milhar
tmp(107) := x"1" & '0' & x"13"; -- LDA @19
tmp(108) := x"8" & '0' & x"0A"; -- CEQ @10      # Compara se o Milhar Ã© igual a 10
tmp(109) := x"7" & '0' & x"71"; -- JEQ @INCREMENTADEZENAMILHAR  # Salta se igual para incrementar a Dezena de Milhar
tmp(110) := x"1" & '0' & x"13"; -- LDA @19
tmp(111) := x"5" & '1' & x"23"; -- STA @291     # Atualiza display HEX3
tmp(112) := x"6" & '0' & x"8F"; -- JMP @RETORNOINCREMENTA
tmp(113) := x"0" & '0' & x"00"; -- NOP #INCREMENTADEZENAMILHAR:pra pular na linha 113
tmp(114) := x"1" & '0' & x"00"; -- LDA @0
tmp(115) := x"5" & '0' & x"13"; -- STA @19      # Reseta o Milhar
tmp(116) := x"5" & '1' & x"23"; -- STA @291     # Atualiza display HEX3
tmp(117) := x"1" & '0' & x"14"; -- LDA @20
tmp(118) := x"2" & '0' & x"01"; -- SOMA @1      # Soma 1 na Dezena de Milhar
tmp(119) := x"5" & '0' & x"14"; -- STA @20      # Armazena o novo valor da Dezena de Milhar
tmp(120) := x"1" & '0' & x"14"; -- LDA @20
tmp(121) := x"8" & '0' & x"0A"; -- CEQ @10      # Compara se a Dezena de Milhar Ã© igual a 10
tmp(122) := x"7" & '0' & x"7E"; -- JEQ @INCREMENTACENTENAMILHAR         # Salta se igual para incrementar a Centena de Milhar
tmp(123) := x"1" & '0' & x"14"; -- LDA @20
tmp(124) := x"5" & '1' & x"24"; -- STA @292     # Atualiza display HEX4
tmp(125) := x"6" & '0' & x"8F"; -- JMP @RETORNOINCREMENTA
tmp(126) := x"0" & '0' & x"00"; -- NOP #INCREMENTACENTENAMILHAR:pra pular na linha 126
tmp(127) := x"1" & '0' & x"00"; -- LDA @0
tmp(128) := x"5" & '0' & x"14"; -- STA @20      # Reseta a Dezena de Milhar
tmp(129) := x"5" & '1' & x"24"; -- STA @292     # Atualiza display HEX4
tmp(130) := x"1" & '0' & x"15"; -- LDA @21
tmp(131) := x"2" & '0' & x"01"; -- SOMA @1      # Soma 1 na Centena de Milhar
tmp(132) := x"5" & '0' & x"15"; -- STA @21      # Armazena o novo valor da Centena de Milhar
tmp(133) := x"1" & '0' & x"15"; -- LDA @21
tmp(134) := x"8" & '0' & x"0A"; -- CEQ @10      # Compara se a Centena de Milhar Ã© igual a 10
tmp(135) := x"7" & '0' & x"8B"; -- JEQ @OVERFLOW        # Salta se igual para tratar overflow
tmp(136) := x"1" & '0' & x"15"; -- LDA @21
tmp(137) := x"5" & '1' & x"25"; -- STA @293     # Atualiza display HEX5
tmp(138) := x"6" & '0' & x"8F"; -- JMP @RETORNOINCREMENTA
tmp(139) := x"0" & '0' & x"00"; -- NOP #OVERFLOW:pra pular na linha 139
tmp(140) := x"1" & '0' & x"01"; -- LDA @1
tmp(141) := x"5" & '1' & x"02"; -- STA @258     # Ativa LEDR9 para indicar overflow
tmp(142) := x"6" & '0' & x"8F"; -- JMP @RETORNOINCREMENTA
tmp(143) := x"0" & '0' & x"00"; -- NOP #RETORNOINCREMENTA:pra pular na linha 143
tmp(144) := x"A" & '0' & x"00"; -- RET
tmp(145) := x"0" & '0' & x"00"; -- NOP #CONFIGURACAO:pra pular na linha 145
tmp(146) := x"1" & '0' & x"00"; -- LDA @0       # Carrega 0
tmp(147) := x"5" & '1' & x"FE"; -- STA @510     # Limpa a leitura de KEY1
tmp(148) := x"5" & '1' & x"20"; -- STA @288     # Limpa display HEX0
tmp(149) := x"5" & '1' & x"21"; -- STA @289     # Limpa display HEX1
tmp(150) := x"5" & '1' & x"22"; -- STA @290     # Limpa display HEX2
tmp(151) := x"5" & '1' & x"23"; -- STA @291     # Limpa display HEX3
tmp(152) := x"5" & '1' & x"24"; -- STA @292     # Limpa display HEX4
tmp(153) := x"5" & '1' & x"25"; -- STA @293     # Limpa display HEX5
tmp(154) := x"0" & '0' & x"00"; -- NOP #AGUARDARKEY1_1:pra pular na linha 154
tmp(155) := x"1" & '1' & x"40"; -- LDA @320     # LÃª o estado dos switches
tmp(156) := x"B" & '0' & x"0F"; -- AND @15      # Aplica mÃ¡scara para isolar os 4 bits inferiores
tmp(157) := x"5" & '0' & x"20"; -- STA @32      # Armazena no endereÃ§o de memÃ³ria dos limites para Unidade
tmp(158) := x"5" & '1' & x"20"; -- STA @288     # Atualiza display HEX0
tmp(159) := x"4" & '0' & x"01"; -- LDI $1
tmp(160) := x"5" & '1' & x"25"; -- STA @293     # Mostra '1' no display HEX5 para indicar configuraÃ§Ã£o da Unidade
tmp(161) := x"1" & '1' & x"61"; -- LDA @353     # LÃª o estado da chave KEY1
tmp(162) := x"8" & '0' & x"01"; -- CEQ @1       # Compara com 1
tmp(163) := x"7" & '0' & x"A5"; -- JEQ @LIMITEDEZ       # Salta se KEY1 pressionado
tmp(164) := x"6" & '0' & x"9A"; -- JMP @AGUARDARKEY1_1
tmp(165) := x"0" & '0' & x"00"; -- NOP #LIMITEDEZ:pra pular na linha 165
tmp(166) := x"1" & '0' & x"00"; -- LDA @0       # Carrega 0
tmp(167) := x"5" & '1' & x"FE"; -- STA @510     # Limpa a leitura de KEY1
tmp(168) := x"0" & '0' & x"00"; -- NOP #AGUARDARKEY1_2:pra pular na linha 168
tmp(169) := x"1" & '1' & x"40"; -- LDA @320     # LÃª o estado dos switches
tmp(170) := x"B" & '0' & x"0F"; -- AND @15      # Aplica mÃ¡scara para isolar os 4 bits inferiores
tmp(171) := x"5" & '0' & x"21"; -- STA @33      # Armazena no endereÃ§o de memÃ³ria dos limites para Dezena
tmp(172) := x"5" & '1' & x"20"; -- STA @288     # Atualiza display HEX0
tmp(173) := x"4" & '0' & x"02"; -- LDI $2
tmp(174) := x"5" & '1' & x"25"; -- STA @293     # Mostra '2' no display HEX5 para indicar configuraÃ§Ã£o da Dezena
tmp(175) := x"1" & '1' & x"61"; -- LDA @353     # LÃª o estado da chave KEY1
tmp(176) := x"8" & '0' & x"01"; -- CEQ @1       # Compara com 1
tmp(177) := x"7" & '0' & x"B3"; -- JEQ @LIMITECEN       # Salta se KEY1 pressionado
tmp(178) := x"6" & '0' & x"A8"; -- JMP @AGUARDARKEY1_2
tmp(179) := x"0" & '0' & x"00"; -- NOP #LIMITECEN:pra pular na linha 179
tmp(180) := x"1" & '0' & x"00"; -- LDA @0       # Carrega 0
tmp(181) := x"5" & '1' & x"FE"; -- STA @510     # Limpa a leitura de KEY1
tmp(182) := x"0" & '0' & x"00"; -- NOP #AGUARDARKEY1_3:pra pular na linha 182
tmp(183) := x"1" & '1' & x"40"; -- LDA @320     # LÃª o estado dos switches
tmp(184) := x"B" & '0' & x"0F"; -- AND @15      # Aplica mÃ¡scara para isolar os 4 bits inferiores
tmp(185) := x"5" & '0' & x"22"; -- STA @34      # Armazena no endereÃ§o de memÃ³ria dos limites para Centena
tmp(186) := x"5" & '1' & x"20"; -- STA @288     # Atualiza display HEX0
tmp(187) := x"4" & '0' & x"03"; -- LDI $3
tmp(188) := x"5" & '1' & x"25"; -- STA @293     # Mostra '3' no display HEX5 para indicar configuraÃ§Ã£o da Centena
tmp(189) := x"1" & '1' & x"61"; -- LDA @353     # LÃª o estado da chave KEY1
tmp(190) := x"8" & '0' & x"01"; -- CEQ @1       # Compara com 1
tmp(191) := x"7" & '0' & x"C1"; -- JEQ @LIMITEUNIM      # Salta se KEY1 pressionado
tmp(192) := x"6" & '0' & x"B6"; -- JMP @AGUARDARKEY1_3
tmp(193) := x"0" & '0' & x"00"; -- NOP #LIMITEUNIM:pra pular na linha 193
tmp(194) := x"1" & '0' & x"00"; -- LDA @0       # Carrega 0
tmp(195) := x"5" & '1' & x"FE"; -- STA @510     # Limpa a leitura de KEY1
tmp(196) := x"0" & '0' & x"00"; -- NOP #AGUARDARKEY1_4:pra pular na linha 196
tmp(197) := x"1" & '1' & x"40"; -- LDA @320     # LÃª o estado dos switches
tmp(198) := x"B" & '0' & x"0F"; -- AND @15      # Aplica mÃ¡scara para isolar os 4 bits inferiores
tmp(199) := x"5" & '0' & x"23"; -- STA @35      # Armazena no endereÃ§o de memÃ³ria dos limites para Unidade de Milhar
tmp(200) := x"5" & '1' & x"20"; -- STA @288     # Atualiza display HEX0
tmp(201) := x"4" & '0' & x"04"; -- LDI $4
tmp(202) := x"5" & '1' & x"25"; -- STA @293     # Mostra '4' no display HEX5 para indicar configuraÃ§Ã£o da Unidade de Milhar
tmp(203) := x"1" & '1' & x"61"; -- LDA @353     # LÃª o estado da chave KEY1
tmp(204) := x"8" & '0' & x"01"; -- CEQ @1       # Compara com 1
tmp(205) := x"7" & '0' & x"CF"; -- JEQ @LIMITEDEZM      # Salta se KEY1 pressionado
tmp(206) := x"6" & '0' & x"C4"; -- JMP @AGUARDARKEY1_4
tmp(207) := x"0" & '0' & x"00"; -- NOP #LIMITEDEZM:pra pular na linha 207
tmp(208) := x"1" & '0' & x"00"; -- LDA @0       # Carrega 0
tmp(209) := x"5" & '1' & x"FE"; -- STA @510     # Limpa a leitura de KEY1
tmp(210) := x"0" & '0' & x"00"; -- NOP #AGUARDARKEY1_5:pra pular na linha 210
tmp(211) := x"1" & '1' & x"40"; -- LDA @320     # LÃª o estado dos switches
tmp(212) := x"B" & '0' & x"0F"; -- AND @15      # Aplica mÃ¡scara para isolar os 4 bits inferiores
tmp(213) := x"5" & '0' & x"24"; -- STA @36      # Armazena no endereÃ§o de memÃ³ria dos limites para Dezena de Milhar
tmp(214) := x"5" & '1' & x"20"; -- STA @288     # Atualiza display HEX0
tmp(215) := x"4" & '0' & x"05"; -- LDI $5
tmp(216) := x"5" & '1' & x"25"; -- STA @293     # Mostra '5' no display HEX5 para indicar configuraÃ§Ã£o da Dezena de Milhar
tmp(217) := x"1" & '1' & x"61"; -- LDA @353     # LÃª o estado da chave KEY1
tmp(218) := x"8" & '0' & x"01"; -- CEQ @1       # Compara com 1
tmp(219) := x"7" & '0' & x"DD"; -- JEQ @LIMITECENM      # Salta se KEY1 pressionado
tmp(220) := x"6" & '0' & x"D2"; -- JMP @AGUARDARKEY1_5
tmp(221) := x"0" & '0' & x"00"; -- NOP #LIMITECENM:pra pular na linha 221
tmp(222) := x"1" & '0' & x"00"; -- LDA @0       # Carrega 0
tmp(223) := x"5" & '1' & x"FE"; -- STA @510     # Limpa a leitura de KEY1
tmp(224) := x"0" & '0' & x"00"; -- NOP #AGUARDARKEY1_6:pra pular na linha 224
tmp(225) := x"1" & '1' & x"40"; -- LDA @320     # LÃª o estado dos switches
tmp(226) := x"B" & '0' & x"0F"; -- AND @15      # Aplica mÃ¡scara para isolar os 4 bits inferiores
tmp(227) := x"5" & '0' & x"25"; -- STA @37      # Armazena no endereÃ§o de memÃ³ria dos limites para Centena de Milhar
tmp(228) := x"5" & '1' & x"20"; -- STA @288     # Atualiza display HEX0
tmp(229) := x"4" & '0' & x"06"; -- LDI $6
tmp(230) := x"5" & '1' & x"25"; -- STA @293     # Mostra '6' no display HEX5 para indicar configuraÃ§Ã£o da Centena de Milhar
tmp(231) := x"1" & '1' & x"61"; -- LDA @353     # LÃª o estado da chave KEY1
tmp(232) := x"8" & '0' & x"01"; -- CEQ @1       # Compara com 1
tmp(233) := x"7" & '0' & x"EB"; -- JEQ @RETORNOCONFIGURACAO     # Salta se KEY1 pressionado
tmp(234) := x"6" & '0' & x"E0"; -- JMP @AGUARDARKEY1_6
tmp(235) := x"0" & '0' & x"00"; -- NOP #RETORNOCONFIGURACAO:pra pular na linha 235
tmp(236) := x"1" & '0' & x"00"; -- LDA @0       # Carrega 0
tmp(237) := x"5" & '1' & x"FE"; -- STA @510     # Limpa a leitura de KEY1
tmp(238) := x"5" & '1' & x"25"; -- STA @293     # Limpa display HEX5
tmp(239) := x"A" & '0' & x"00"; -- RET
tmp(240) := x"0" & '0' & x"00"; -- NOP #REINICIACONTAGEM:pra pular na linha 240
tmp(241) := x"1" & '0' & x"00"; -- LDA @0
tmp(242) := x"5" & '1' & x"FD"; -- STA @509     # Limpa valor no endereÃ§o 509
tmp(243) := x"5" & '0' & x"10"; -- STA @16      # Reseta contador de Unidade
tmp(244) := x"5" & '0' & x"11"; -- STA @17      # Reseta contador de Dezena
tmp(245) := x"5" & '0' & x"12"; -- STA @18      # Reseta contador de Centena
tmp(246) := x"5" & '0' & x"13"; -- STA @19      # Reseta contador de Milhar
tmp(247) := x"5" & '0' & x"14"; -- STA @20      # Reseta contador de Dezena de Milhar
tmp(248) := x"5" & '0' & x"15"; -- STA @21      # Reseta contador de Centena de Milhar
tmp(249) := x"5" & '1' & x"20"; -- STA @288     # Limpa display HEX0
tmp(250) := x"5" & '1' & x"21"; -- STA @289     # Limpa display HEX1
tmp(251) := x"5" & '1' & x"22"; -- STA @290     # Limpa display HEX2
tmp(252) := x"5" & '1' & x"23"; -- STA @291     # Limpa display HEX3
tmp(253) := x"5" & '1' & x"24"; -- STA @292     # Limpa display HEX4
tmp(254) := x"5" & '1' & x"25"; -- STA @293     # Limpa display HEX5
tmp(255) := x"5" & '0' & x"1B"; -- STA @27      # Limpa a flag de limite
tmp(256) := x"5" & '1' & x"01"; -- STA @257     # Limpa LEDR8
tmp(257) := x"5" & '1' & x"02"; -- STA @258     # Limpa LEDR9
tmp(258) := x"A" & '0' & x"00"; -- RET
tmp(259) := x"0" & '0' & x"00"; -- NOP #VERIFICARLIMITE:pra pular na linha 259
tmp(260) := x"1" & '0' & x"10"; -- LDA @16      # Carrega valor da Unidade
tmp(261) := x"8" & '0' & x"20"; -- CEQ @32      # Compara com o limite para Unidade
tmp(262) := x"7" & '1' & x"08"; -- JEQ @VERDEZENAS      # Salta se igual para verificar limite de Dezena
tmp(263) := x"6" & '1' & x"25"; -- JMP @RETORNOVERIFICALIMITE
tmp(264) := x"0" & '0' & x"00"; -- NOP #VERDEZENAS:pra pular na linha 264
tmp(265) := x"1" & '0' & x"11"; -- LDA @17      # Carrega valor da Dezena
tmp(266) := x"8" & '0' & x"21"; -- CEQ @33      # Compara com o limite para Dezena
tmp(267) := x"7" & '1' & x"0D"; -- JEQ @VERCENTENAS     # Salta se igual para verificar limite de Centena
tmp(268) := x"6" & '1' & x"25"; -- JMP @RETORNOVERIFICALIMITE
tmp(269) := x"0" & '0' & x"00"; -- NOP #VERCENTENAS:pra pular na linha 269
tmp(270) := x"1" & '0' & x"12"; -- LDA @18      # Carrega valor da Centena
tmp(271) := x"8" & '0' & x"22"; -- CEQ @34      # Compara com o limite para Centena
tmp(272) := x"7" & '1' & x"12"; -- JEQ @VERUNIDADESM    # Salta se igual para verificar limite de Unidade de Milhar
tmp(273) := x"6" & '1' & x"25"; -- JMP @RETORNOVERIFICALIMITE
tmp(274) := x"0" & '0' & x"00"; -- NOP #VERUNIDADESM:pra pular na linha 274
tmp(275) := x"1" & '0' & x"13"; -- LDA @19      # Carrega valor da Unidade de Milhar
tmp(276) := x"8" & '0' & x"23"; -- CEQ @35      # Compara com o limite para Unidade de Milhar
tmp(277) := x"7" & '1' & x"17"; -- JEQ @VERDEZENASM     # Salta se igual para verificar limite de Dezena de Milhar
tmp(278) := x"6" & '1' & x"25"; -- JMP @RETORNOVERIFICALIMITE
tmp(279) := x"0" & '0' & x"00"; -- NOP #VERDEZENASM:pra pular na linha 279
tmp(280) := x"1" & '0' & x"14"; -- LDA @20      # Carrega valor da Dezena de Milhar
tmp(281) := x"8" & '0' & x"24"; -- CEQ @36      # Compara com o limite para Dezena de Milhar
tmp(282) := x"7" & '1' & x"1C"; -- JEQ @VERCENTENASM    # Salta se igual para verificar limite de Centena de Milhar
tmp(283) := x"6" & '1' & x"25"; -- JMP @RETORNOVERIFICALIMITE
tmp(284) := x"0" & '0' & x"00"; -- NOP #VERCENTENASM:pra pular na linha 284
tmp(285) := x"1" & '0' & x"15"; -- LDA @21      # Carrega valor da Centena de Milhar
tmp(286) := x"8" & '0' & x"25"; -- CEQ @37      # Compara com o limite para Centena de Milhar
tmp(287) := x"7" & '1' & x"21"; -- JEQ @LIGARFLAG       # Salta se igual para ativar flag de limite
tmp(288) := x"6" & '1' & x"25"; -- JMP @RETORNOVERIFICALIMITE
tmp(289) := x"0" & '0' & x"00"; -- NOP #LIGARFLAG:pra pular na linha 289
tmp(290) := x"1" & '0' & x"01"; -- LDA @1
tmp(291) := x"5" & '0' & x"1B"; -- STA @27      # Ativa a flag de limite
tmp(292) := x"5" & '1' & x"01"; -- STA @257     # Ativa LEDR8 para indicar o limite atingido
tmp(293) := x"0" & '0' & x"00"; -- NOP #RETORNOVERIFICALIMITE:pra pular na linha 293
tmp(294) := x"A" & '0' & x"00"; -- RET
	return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;